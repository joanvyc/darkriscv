/*
 * Copyright (c) 2018, Marcelo Samsoniuk
 * All rights reserved.
 * 
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions are met:
 * 
 * * Redistributions of source code must retain the above copyright notice, this
 *   list of conditions and the following disclaimer.
 * 
 * * Redistributions in binary form must reproduce the above copyright notice,
 *   this list of conditions and the following disclaimer in the documentation
 *   and/or other materials provided with the distribution.
 * 
 * * Neither the name of the copyright holder nor the names of its
 *   contributors may be used to endorse or promote products derived from
 *   this software without specific prior written permission.
 * 
 * THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 * AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 * DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 * FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 * DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 * SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 * CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 * OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 * OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE. 
 */

`timescale 1ns / 1ps

// implemented opcodes:

`define LUI     7'b01101_11      // lui   rd,imm[31:12]
`define AUIPC   7'b00101_11      // auipc rd,imm[31:12]
`define JAL     7'b11011_11      // jal   rd,imm[xxxxx]
`define JALR    7'b11001_11      // jalr  rd,rs1,imm[11:0] 
`define BCC     7'b11000_11      // bcc   rs1,rs2,imm[12:1]
`define LCC     7'b00000_11      // lxx   rd,rs1,imm[11:0]
`define SCC     7'b01000_11      // sxx   rs1,rs2,imm[11:0]
`define MCC     7'b00100_11      // xxxi  rd,rs1,imm[11:0]
`define RCC     7'b01100_11      // xxx   rd,rs1,rs2 
`define MAC     7'b11111_11      // mac   rd,rs1,rs2

// not implemented opcodes:

`define FCC     7'b00011_11      // fencex
`define CCC     7'b11100_11      // exx, csrxx

// configuration file

`include "config.vh"

module darkfetch
//#(
//    parameter [31:0] RESET_PC = 0,
//    parameter [31:0] RESET_SP = 4096
//) 
(
    input             clk,   // clock
    input             res,   // reset

	input             en,
	output			  valid,
	
	darkbus.prov	  bus,
	
	// Instruction data (in)
	input 			  pc,
	
	// Instruction data (out)
	output			  pc_o,
	output 		      inst
);

	typedef enum logic [1:0] {IDLE, EXEC} fetch_state;
	
	fetch_state  curr_st, next_st;

	logic [31:0] curr_pc, next_pc;
	logic [31:0] curr_inst, next_inst;	
	
	assign bus.data = 32'bZ;
	
	assign pc_o = curr_pc;
	assign inst = curr_inst;
	
	always_comb
	begin
		case (curr_st) 
			IDLE:
				begin
					if (en) begin
						next_pc = pc;
						next_st = EXEC;
						next_inst = curr_inst;
					end	else begin
						next_pc = curr_pc;
						next_st = curr_st;
						next_inst = curr_inst;
					end
                end
			default: 
				begin
					if (bus.valid) begin
						next_pc = curr_pc;
						next_st = IDLE;
						next_inst = bus.data;
					end else begin
						next_pc = curr_pc;
						next_st = curr_st;
						next_inst = curr_inst;
					end
				end
		endcase
	end
	
	always @(posedge clk)
	begin
		curr_pc <= next_pc;
		curr_st <= next_st;
		curr_inst <= next_inst;
	end
	
	always_comb
	begin
		case (curr_st)
			IDLE:
				begin
					bus.en = 0;
					bus.rw = 0;
				end
			default:
				begin
					bus.en = 1;
					bus.rw = 0;
					bus.addr = curr_pc;
				end
		endcase
	end
	
endmodule
