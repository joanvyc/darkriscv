/*
 * Copyright (c) 2021, Joan Vinyals Ylla-Catala
 * All rights reserved.
 * 
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions are met:
 * 
 * * Redistributions of source code must retain the above copyright notice, this
 *   list of conditions and the following disclaimer.
 * 
 * * Redistributions in binary form must reproduce the above copyright notice,
 *   this list of conditions and the following disclaimer in the documentation
 *   and/or other materials provided with the distribution.
 * 
 * * Neither the name of the copyright holder nor the names of its
 *   contributors may be used to endorse or promote products derived from
 *   this software without specific prior written permission.
 * 
 * THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 * AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
 * DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
 * FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 * DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
 * SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
 * CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 * OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
 * OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE. 
 */

module darkocrom
(
  input           XCLK,
  input           XRES,

  input           EN,
  input           RD,
  input           WR,

  input  [3:0]    BE,

  output          ACK,

  input  [31:0]   addr,
  inout  [31:0]   data

`ifdef _EXTERNAL_RAM_
  ,darkaxi.Master  ram
`endif

);

`ifdef _EXTERNAL_RAM_


`else

  (* ram_style = "block" *) reg [31:0] MEM [0:511];

  assign data = (EN && RD) ? MEM[addr[31:2]] : 32'bz;

  always @(posedge XCLK)
  begin
    if (EN && WE)
    begin
      if (BE)
      begin
        integer i;
        for (i=0; i!=4; i=i+1)
        begin
          if (BE[i]) MEM[addr[31:2]][i * 8 + 7: i * 8] = data[i * 8 + 7: i * 8];
        end
      end

      else
        MEM[addr[31:2]] = data;
    end
  end

`endif

endmodule
